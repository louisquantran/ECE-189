`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/31/2025 03:30:11 PM
// Design Name: 
// Module Name: Fetch
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Fetch(
    input logic clk,
    input logic reset,
    
    // Downstream    
    input logic [31:0] PC_in,
    
    // Upstream
    input logic ready_in,
    output logic [31:0] instr_out,
    output logic [31:0] PC_out,
    output logic [31:0] PC_4,
    output logic valid_out,
);
    logic [31:0] PC_buf;
    logic [31:0] instr_buf;
    logic valid_out_buf;
    logic [31:0] PC_icache;
    logic [31:0] instr_icache;
    
    // Call ICache
    ICache ICache_dut (
        .clk(clk),
        .reset(reset),
        .address(PC_in),
        .instruction(instr_icache)
    );
    
    // Combinational assignments
    assign PC_out = PC_buf;
    assign PC_4 = PC_buf + 32'd4;
    assign valid_out = valid_out_buf;
    assign instr_out = instr_buf;
    
    // Sequential assignments
    always_ff @(posedge clk) begin
        if (reset) begin
            valid_out_buf <= 1'b0;  
            instr_buf <= 32'b0;
            PC_buf <= 32'b0;
        end else begin
            PC_icache <= PC_in;
            if (!valid_out_buf || ready_in) begin
                valid_out_buf <= 1'b1;
                PC_buf <= PC_icache;
                instr_buf <= instr_icache;
            end
        end
    end
endmodule